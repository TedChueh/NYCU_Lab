module bit_invert (
    input in0,
    output out0
);

not g1(out0, in0);
    
endmodule